`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Gunnar Pederson
// 
// Create Date: 05/28/2021 11:54:53 AM
// Design Name: 
// Module Name: mux_8_1
// Project Name: project 5 Mux Demux circuit
// Target Devices: 
// Tool Versions: Vivado 2020.2
// Description: mux 8 to 1
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_8_1(
    input [7:0] I,      //input
    input [2:0] S,      //mux select
    output Y            //mux output
    );
    
reg tmp;
    
always @ (S, I)
begin
    case (S)
    3'b000: tmp <= I[0];
    3'b001: tmp <= I[1];
    3'b010: tmp <= I[2];
    3'b011: tmp <= I[3];
    3'b100: tmp <= I[4];
    3'b101: tmp <= I[5];
    3'b110: tmp <= I[6];
    3'b111: tmp <= I[7];
    default: tmp <= 0;
    endcase
end 
    
assign Y = tmp;
    
endmodule
